--
-- VHDL Architecture OBC_test.test.SPI_tester
--
-- Created:
--          by - Lucas.Mayor (DESKTOP-3I0F3HP)
--          at - 13:14:41 13.07.2020
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE SPI_tester OF test IS
BEGIN
END ARCHITECTURE SPI_tester;

